library verilog;
use verilog.vl_types.all;
entity nol_11011_mealy is
end nol_11011_mealy;
