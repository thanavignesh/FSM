library verilog;
use verilog.vl_types.all;
entity ol_11011_mealy is
end ol_11011_mealy;
