library verilog;
use verilog.vl_types.all;
entity nol_1101_moore is
end nol_1101_moore;
