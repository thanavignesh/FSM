library verilog;
use verilog.vl_types.all;
entity ol_11011_moore is
end ol_11011_moore;
