library verilog;
use verilog.vl_types.all;
entity nol_1101_mealy is
end nol_1101_mealy;
