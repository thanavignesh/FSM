library verilog;
use verilog.vl_types.all;
entity ol_1101_moore is
end ol_1101_moore;
