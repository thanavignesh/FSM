library verilog;
use verilog.vl_types.all;
entity mealy_fsm_tb is
end mealy_fsm_tb;
