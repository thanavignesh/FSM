library verilog;
use verilog.vl_types.all;
entity moore_tb is
end moore_tb;
