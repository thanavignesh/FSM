library verilog;
use verilog.vl_types.all;
entity nol_11011_moore is
end nol_11011_moore;
